module test (o, x, y);
    output o;
    input x, y;

    and a1 (o, x ,y);
endmodule
